// megafunction wizard: %ALTSQRT%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altsqrt 

// ============================================================
// File Name: Sqrt_64b.v
// Megafunction Name(s):
// 			altsqrt
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 7.2 Build 151 09/26/2007 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2007 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module Sqrt_64b (
	clk,
	radical,
	q,
	remainder);

	input	  clk;
	input	[63:0]  radical;
	output	[31:0]  q;
	output	[32:0]  remainder;

	wire [32:0] sub_wire0;
	wire [31:0] sub_wire1;
	wire [32:0] remainder = sub_wire0[32:0];
	wire [31:0] q = sub_wire1[31:0];

	altsqrt	altsqrt_component (
				.radical (radical),
				.clk (clk),
				.remainder (sub_wire0),
				.q (sub_wire1)
				// synopsys translate_off
				,
				.aclr (),
				.ena ()
				// synopsys translate_on
				);
	defparam
		altsqrt_component.pipeline = 10,
		altsqrt_component.q_port_width = 32,
		altsqrt_component.r_port_width = 33,
		altsqrt_component.width = 64;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix II"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "1"
// Retrieval info: CONSTANT: PIPELINE NUMERIC "10"
// Retrieval info: CONSTANT: Q_PORT_WIDTH NUMERIC "32"
// Retrieval info: CONSTANT: R_PORT_WIDTH NUMERIC "33"
// Retrieval info: CONSTANT: WIDTH NUMERIC "64"
// Retrieval info: USED_PORT: clk 0 0 0 0 INPUT NODEFVAL clk
// Retrieval info: USED_PORT: q 0 0 32 0 OUTPUT NODEFVAL q[31..0]
// Retrieval info: USED_PORT: radical 0 0 64 0 INPUT NODEFVAL radical[63..0]
// Retrieval info: USED_PORT: remainder 0 0 33 0 OUTPUT NODEFVAL remainder[32..0]
// Retrieval info: CONNECT: @clk 0 0 0 0 clk 0 0 0 0
// Retrieval info: CONNECT: @radical 0 0 64 0 radical 0 0 64 0
// Retrieval info: CONNECT: q 0 0 32 0 @q 0 0 32 0
// Retrieval info: CONNECT: remainder 0 0 33 0 @remainder 0 0 33 0
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL Sqrt_64b.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL Sqrt_64b.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Sqrt_64b.cmp TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL Sqrt_64b.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Sqrt_64b_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Sqrt_64b_bb.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL Sqrt_64b_syn.v TRUE
// Retrieval info: LIB_FILE: altera_mf
